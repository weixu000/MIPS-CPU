module ROM(
    input [30:0] addr,
    output [31:0] data
);

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [ROM_SIZE:0] ROMDATA[ROM_SIZE-1:0];

assign data = addr[30:2]<ROM_SIZE ? ROMDATA[addr[30:2]] : 32'b0;

integer i;
initial begin
    ROMDATA[0] <= 32'h08000002;
    ROMDATA[1] <= 32'h0800001f;
    ROMDATA[2] <= 32'h3c084000;
    ROMDATA[3] <= 32'h2109000c;
    ROMDATA[4] <= 32'h210a001a;
    ROMDATA[5] <= 32'h210b0018;
    ROMDATA[6] <= 32'h210c001c;
    ROMDATA[7] <= 32'h200d0000;
    ROMDATA[8] <= 32'h3c0effff;
    ROMDATA[9] <= 32'h35ce3caf;
    ROMDATA[10] <= 32'had0e0000;
    ROMDATA[11] <= 32'h3c0effff;
    ROMDATA[12] <= 32'h35ceffff;
    ROMDATA[13] <= 32'had0e0004;
    ROMDATA[14] <= 32'h200e0003;
    ROMDATA[15] <= 32'had0e0008;
    ROMDATA[16] <= 32'h201f004c;
    ROMDATA[17] <= 32'had0e0008;
    ROMDATA[18] <= 32'h03e00008;
    ROMDATA[19] <= 32'h8d0e0020;
    ROMDATA[20] <= 32'h000e70c2;
    ROMDATA[21] <= 32'h21ceffff;
    ROMDATA[22] <= 32'h11c00001;
    ROMDATA[23] <= 32'h08000013;
    ROMDATA[24] <= 32'h11a00003;
    ROMDATA[25] <= 32'h200d0000;
    ROMDATA[26] <= 32'h8d910000;
    ROMDATA[27] <= 32'h0800007f;
    ROMDATA[28] <= 32'h8d900000;
    ROMDATA[29] <= 32'h21ad0001;
    ROMDATA[30] <= 32'h08000013;
    ROMDATA[31] <= 32'h200e0000;
    ROMDATA[32] <= 32'had0e0008;
    ROMDATA[33] <= 32'h11a00006;
    ROMDATA[34] <= 32'h21aeffff;
    ROMDATA[35] <= 32'h11c0000e;
    ROMDATA[36] <= 32'h21aefffe;
    ROMDATA[37] <= 32'h11c00015;
    ROMDATA[38] <= 32'h21aefffd;
    ROMDATA[39] <= 32'h11c0001d;
    ROMDATA[40] <= 32'h00109700;
    ROMDATA[41] <= 32'h00129702;
    ROMDATA[42] <= 32'h0c00004e;
    ROMDATA[43] <= 32'h22520e00;
    ROMDATA[44] <= 32'had520000;
    ROMDATA[45] <= 32'h21ad0001;
    ROMDATA[46] <= 32'h200e0003;
    ROMDATA[47] <= 32'had0e0008;
    ROMDATA[48] <= 32'h235afffc;
    ROMDATA[49] <= 32'h03400008;
    ROMDATA[50] <= 32'h00109102;
    ROMDATA[51] <= 32'h0c00004e;
    ROMDATA[52] <= 32'h22520d00;
    ROMDATA[53] <= 32'had520000;
    ROMDATA[54] <= 32'h21ad0001;
    ROMDATA[55] <= 32'h200e0003;
    ROMDATA[56] <= 32'had0e0008;
    ROMDATA[57] <= 32'h235afffc;
    ROMDATA[58] <= 32'h03400008;
    ROMDATA[59] <= 32'h00119700;
    ROMDATA[60] <= 32'h00129702;
    ROMDATA[61] <= 32'h0c00004e;
    ROMDATA[62] <= 32'h22520b00;
    ROMDATA[63] <= 32'had520000;
    ROMDATA[64] <= 32'h21ad0001;
    ROMDATA[65] <= 32'h200e0003;
    ROMDATA[66] <= 32'had0e0008;
    ROMDATA[67] <= 32'h235afffc;
    ROMDATA[68] <= 32'h03400008;
    ROMDATA[69] <= 32'h00119102;
    ROMDATA[70] <= 32'h0c00004e;
    ROMDATA[71] <= 32'h22520700;
    ROMDATA[72] <= 32'had520000;
    ROMDATA[73] <= 32'h200d0000;
    ROMDATA[74] <= 32'h200e0003;
    ROMDATA[75] <= 32'had0e0008;
    ROMDATA[76] <= 32'h235afffc;
    ROMDATA[77] <= 32'h03400008;
    ROMDATA[78] <= 32'h200f0002;
    ROMDATA[79] <= 32'h1240002d;
    ROMDATA[80] <= 32'h200f009e;
    ROMDATA[81] <= 32'h2258ffff;
    ROMDATA[82] <= 32'h1300002a;
    ROMDATA[83] <= 32'h200f0024;
    ROMDATA[84] <= 32'h2258fffe;
    ROMDATA[85] <= 32'h13000027;
    ROMDATA[86] <= 32'h200f000c;
    ROMDATA[87] <= 32'h2258fffd;
    ROMDATA[88] <= 32'h13000024;
    ROMDATA[89] <= 32'h200f0098;
    ROMDATA[90] <= 32'h2258fffc;
    ROMDATA[91] <= 32'h13000021;
    ROMDATA[92] <= 32'h200f0048;
    ROMDATA[93] <= 32'h2258fffb;
    ROMDATA[94] <= 32'h1300001e;
    ROMDATA[95] <= 32'h200f0040;
    ROMDATA[96] <= 32'h2258fffa;
    ROMDATA[97] <= 32'h1300001b;
    ROMDATA[98] <= 32'h200f001e;
    ROMDATA[99] <= 32'h2258fff9;
    ROMDATA[100] <= 32'h13000018;
    ROMDATA[101] <= 32'h200f0000;
    ROMDATA[102] <= 32'h2258fff8;
    ROMDATA[103] <= 32'h13000015;
    ROMDATA[104] <= 32'h200f0004;
    ROMDATA[105] <= 32'h2258fff7;
    ROMDATA[106] <= 32'h13000012;
    ROMDATA[107] <= 32'h200f0008;
    ROMDATA[108] <= 32'h2258fff6;
    ROMDATA[109] <= 32'h1300000f;
    ROMDATA[110] <= 32'h200f00c0;
    ROMDATA[111] <= 32'h2258fff5;
    ROMDATA[112] <= 32'h1300000c;
    ROMDATA[113] <= 32'h200f0062;
    ROMDATA[114] <= 32'h2258fff4;
    ROMDATA[115] <= 32'h13000009;
    ROMDATA[116] <= 32'h200f0084;
    ROMDATA[117] <= 32'h2258fff3;
    ROMDATA[118] <= 32'h13000006;
    ROMDATA[119] <= 32'h200f0062;
    ROMDATA[120] <= 32'h2258fff2;
    ROMDATA[121] <= 32'h13000003;
    ROMDATA[122] <= 32'h200f0072;
    ROMDATA[123] <= 32'h2258fff1;
    ROMDATA[124] <= 32'h13000000;
    ROMDATA[125] <= 32'h000f9020;
    ROMDATA[126] <= 32'h03e00008;
    ROMDATA[127] <= 32'h12110009;
    ROMDATA[128] <= 32'h1e110004;
    ROMDATA[129] <= 32'h02307822;
    ROMDATA[130] <= 32'h120f0008;
    ROMDATA[131] <= 32'h21f10000;
    ROMDATA[132] <= 32'h08000080;
    ROMDATA[133] <= 32'h02117822;
    ROMDATA[134] <= 32'h122f0004;
    ROMDATA[135] <= 32'h21f00000;
    ROMDATA[136] <= 32'h08000080;
    ROMDATA[137] <= 32'h22040000;
    ROMDATA[138] <= 32'h208f0000;
    ROMDATA[139] <= 32'h21e40000;
    ROMDATA[140] <= 32'had240000;
    ROMDATA[141] <= 32'had640000;
    ROMDATA[142] <= 32'h1000ffff;
    for (i=143; i<ROM_SIZE; i=i+1) begin
        ROMDATA[i] <= 32'b0;
    end
end
endmodule
