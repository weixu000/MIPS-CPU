module ROM(
    input [30:0] addr,
    output [31:0] data
);

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data = addr[30:2]<ROM_SIZE ? ROMDATA[addr[30:2]] : 32'b0;

integer i;
initial begin
    ROMDATA[0] <= 32'h08000002;
    ROMDATA[1] <= 32'h0800001f;
    ROMDATA[2] <= 32'h3c084000;
    ROMDATA[3] <= 32'h2109000c;
    ROMDATA[4] <= 32'h210a0014;
    ROMDATA[5] <= 32'h210c001c;
    ROMDATA[6] <= 32'h200d0000;
    ROMDATA[7] <= 32'h20190000;
    ROMDATA[8] <= 32'h3c0effff;
    ROMDATA[9] <= 32'h35ce3caf;
    ROMDATA[10] <= 32'had0e0000;
    ROMDATA[11] <= 32'h3c0effff;
    ROMDATA[12] <= 32'h35ceffff;
    ROMDATA[13] <= 32'had0e0004;
    ROMDATA[14] <= 32'h200e0003;
    ROMDATA[15] <= 32'had0e0008;
    ROMDATA[16] <= 32'h201f004c;
    ROMDATA[17] <= 32'had0e0008;
    ROMDATA[18] <= 32'h03e00008;
    ROMDATA[19] <= 32'h8d0e0020;
    ROMDATA[20] <= 32'h000e70c2;
    ROMDATA[21] <= 32'h21ceffff;
    ROMDATA[22] <= 32'h00000000;
    ROMDATA[23] <= 32'h11c00001;
    ROMDATA[24] <= 32'h08000013;
    ROMDATA[25] <= 32'h13200002;
    ROMDATA[26] <= 32'h8d910000;
    ROMDATA[27] <= 32'h08000095;
    ROMDATA[28] <= 32'h8d900000;
    ROMDATA[29] <= 32'h23390001;
    ROMDATA[30] <= 32'h08000013;
    ROMDATA[31] <= 32'h200e0000;
    ROMDATA[32] <= 32'had0e0008;
    ROMDATA[33] <= 32'h11a00009;
    ROMDATA[34] <= 32'h21aeffff;
    ROMDATA[35] <= 32'h00000000;
    ROMDATA[36] <= 32'h11c00011;
    ROMDATA[37] <= 32'h21aefffe;
    ROMDATA[38] <= 32'h00000000;
    ROMDATA[39] <= 32'h11c00018;
    ROMDATA[40] <= 32'h21aefffd;
    ROMDATA[41] <= 32'h00000000;
    ROMDATA[42] <= 32'h11c00020;
    ROMDATA[43] <= 32'h00109700;
    ROMDATA[44] <= 32'h00129702;
    ROMDATA[45] <= 32'h0c000055;
    ROMDATA[46] <= 32'h22520e00;
    ROMDATA[47] <= 32'had520000;
    ROMDATA[48] <= 32'h21ad0001;
    ROMDATA[49] <= 32'h200e0003;
    ROMDATA[50] <= 32'had0e0008;
    ROMDATA[51] <= 32'h235afffc;
    ROMDATA[52] <= 32'h00000000;
    ROMDATA[53] <= 32'h03400008;
    ROMDATA[54] <= 32'h00109102;
    ROMDATA[55] <= 32'h0c000055;
    ROMDATA[56] <= 32'h22520d00;
    ROMDATA[57] <= 32'had520000;
    ROMDATA[58] <= 32'h21ad0001;
    ROMDATA[59] <= 32'h200e0003;
    ROMDATA[60] <= 32'had0e0008;
    ROMDATA[61] <= 32'h235afffc;
    ROMDATA[62] <= 32'h00000000;
    ROMDATA[63] <= 32'h03400008;
    ROMDATA[64] <= 32'h00119700;
    ROMDATA[65] <= 32'h00129702;
    ROMDATA[66] <= 32'h0c000055;
    ROMDATA[67] <= 32'h22520b00;
    ROMDATA[68] <= 32'had520000;
    ROMDATA[69] <= 32'h21ad0001;
    ROMDATA[70] <= 32'h200e0003;
    ROMDATA[71] <= 32'had0e0008;
    ROMDATA[72] <= 32'h235afffc;
    ROMDATA[73] <= 32'h00000000;
    ROMDATA[74] <= 32'h03400008;
    ROMDATA[75] <= 32'h00119102;
    ROMDATA[76] <= 32'h0c000055;
    ROMDATA[77] <= 32'h22520700;
    ROMDATA[78] <= 32'had520000;
    ROMDATA[79] <= 32'h200d0000;
    ROMDATA[80] <= 32'h200e0003;
    ROMDATA[81] <= 32'had0e0008;
    ROMDATA[82] <= 32'h235afffc;
    ROMDATA[83] <= 32'h00000000;
    ROMDATA[84] <= 32'h03400008;
    ROMDATA[85] <= 32'h200f0003;
    ROMDATA[86] <= 32'h1240003c;
    ROMDATA[87] <= 32'h200f009f;
    ROMDATA[88] <= 32'h2258ffff;
    ROMDATA[89] <= 32'h00000000;
    ROMDATA[90] <= 32'h13000038;
    ROMDATA[91] <= 32'h200f0025;
    ROMDATA[92] <= 32'h2258fffe;
    ROMDATA[93] <= 32'h00000000;
    ROMDATA[94] <= 32'h13000034;
    ROMDATA[95] <= 32'h200f000d;
    ROMDATA[96] <= 32'h2258fffd;
    ROMDATA[97] <= 32'h00000000;
    ROMDATA[98] <= 32'h13000030;
    ROMDATA[99] <= 32'h200f0099;
    ROMDATA[100] <= 32'h2258fffc;
    ROMDATA[101] <= 32'h00000000;
    ROMDATA[102] <= 32'h1300002c;
    ROMDATA[103] <= 32'h200f0049;
    ROMDATA[104] <= 32'h2258fffb;
    ROMDATA[105] <= 32'h00000000;
    ROMDATA[106] <= 32'h13000028;
    ROMDATA[107] <= 32'h200f0041;
    ROMDATA[108] <= 32'h2258fffa;
    ROMDATA[109] <= 32'h00000000;
    ROMDATA[110] <= 32'h13000024;
    ROMDATA[111] <= 32'h200f001f;
    ROMDATA[112] <= 32'h2258fff9;
    ROMDATA[113] <= 32'h00000000;
    ROMDATA[114] <= 32'h13000020;
    ROMDATA[115] <= 32'h200f0001;
    ROMDATA[116] <= 32'h2258fff8;
    ROMDATA[117] <= 32'h00000000;
    ROMDATA[118] <= 32'h1300001c;
    ROMDATA[119] <= 32'h200f0009;
    ROMDATA[120] <= 32'h2258fff7;
    ROMDATA[121] <= 32'h00000000;
    ROMDATA[122] <= 32'h13000018;
    ROMDATA[123] <= 32'h200f0011;
    ROMDATA[124] <= 32'h2258fff6;
    ROMDATA[125] <= 32'h00000000;
    ROMDATA[126] <= 32'h13000014;
    ROMDATA[127] <= 32'h200f00c1;
    ROMDATA[128] <= 32'h2258fff5;
    ROMDATA[129] <= 32'h00000000;
    ROMDATA[130] <= 32'h13000010;
    ROMDATA[131] <= 32'h200f0063;
    ROMDATA[132] <= 32'h2258fff4;
    ROMDATA[133] <= 32'h00000000;
    ROMDATA[134] <= 32'h1300000c;
    ROMDATA[135] <= 32'h200f0085;
    ROMDATA[136] <= 32'h2258fff3;
    ROMDATA[137] <= 32'h00000000;
    ROMDATA[138] <= 32'h13000008;
    ROMDATA[139] <= 32'h200f0061;
    ROMDATA[140] <= 32'h2258fff2;
    ROMDATA[141] <= 32'h00000000;
    ROMDATA[142] <= 32'h13000004;
    ROMDATA[143] <= 32'h200f0071;
    ROMDATA[144] <= 32'h2258fff1;
    ROMDATA[145] <= 32'h00000000;
    ROMDATA[146] <= 32'h13000000;
    ROMDATA[147] <= 32'h000f9020;
    ROMDATA[148] <= 32'h03e00008;
    ROMDATA[149] <= 32'h1211000e;
    ROMDATA[150] <= 32'h22130000;
    ROMDATA[151] <= 32'h22340000;
    ROMDATA[152] <= 32'h00000000;
    ROMDATA[153] <= 32'h1e740005;
    ROMDATA[154] <= 32'h02935822;
    ROMDATA[155] <= 32'h00000000;
    ROMDATA[156] <= 32'h126b0009;
    ROMDATA[157] <= 32'h21740000;
    ROMDATA[158] <= 32'h08000098;
    ROMDATA[159] <= 32'h02745822;
    ROMDATA[160] <= 32'h00000000;
    ROMDATA[161] <= 32'h128b0004;
    ROMDATA[162] <= 32'h21730000;
    ROMDATA[163] <= 32'h08000098;
    ROMDATA[164] <= 32'h22240000;
    ROMDATA[165] <= 32'h208b0000;
    ROMDATA[166] <= 32'h21640000;
    ROMDATA[167] <= 32'had240000;
    ROMDATA[168] <= 32'had040018;
    ROMDATA[169] <= 32'h20000000;
    ROMDATA[170] <= 32'h1000fffe;
    for (i=171; i<ROM_SIZE; i=i+1) begin
        ROMDATA[i] <= 32'b0;
    end
end
endmodule
